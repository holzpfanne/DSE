-------------------------------------------------------------------------------
--                                                                      
--                        JK Flip flop
--  
-------------------------------------------------------------------------------

configuration JK_struc_cfg of JK is
  for struc        -- architecture struc is used for entity data_bus
  end for;
end JK_struc_cfg;

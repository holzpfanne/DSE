-------------------------------------------------------------------------------
--                                                                      
--                        JK and D Flip flop
--  
-------------------------------------------------------------------------------

configuration four_struc_cfg of four is
  for struc        
  end for;
end four_struc_cfg;

-------------------------------------------------------------------------------
--                                                                      
--                        D Flip flop
--  
-------------------------------------------------------------------------------

configuration D_struc_cfg of D is
  for struc        
  end for;
end D_struc_cfg;

-------------------------------------------------------------------------------
--                                                                      
--                        calucator project
--  
-------------------------------------------------------------------------------

configuration calc_rtl_cfg of io_ctrl is
  for rtl        -- architecture rtl is used for entity data_bus
  end for;
end calc_rtl_cfg;

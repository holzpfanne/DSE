-------------------------------------------------------------------------------
--                                                                      
--                        8-bit Adder
--  
-------------------------------------------------------------------------------

configuration eight_bit_struc_cfg of eight_bit is
  for struc        
  end for;
end eight_bit_struc_cfg;

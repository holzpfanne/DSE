-------------------------------------------------------------------------------
--                                                                      
--                        calucator project
--  
-------------------------------------------------------------------------------

configuration calculator_rtl_cfg of calculator is
  for rtl        -- architecture rtl is used for entity data_bus
  end for;
end calculator_rtl_cfg;

-------------------------------------------------------------------------------
--                                                                      
--                        calucator project
--  
-------------------------------------------------------------------------------

configuration calc_rtl_cfg of calc is
  for rtl        -- architecture rtl is used for entity data_bus
  end for;
end calc_rtl_cfg;

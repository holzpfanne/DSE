-------------------------------------------------------------------------------
--                                                                      
--                        JK and D Flip flop
--  
-------------------------------------------------------------------------------

configuration JKD_struc_cfg of JKD is
  for struc        
  end for;
end JKD_struc_cfg;

-------------------------------------------------------------------------------
--                                                                      
--                        ocalucator project, calc_ctrl
--  
-------------------------------------------------------------------------------

configuration calc_ctrl_rtl_cfg of calc_ctrl is
  for rtl        -- architecture rtl is used for entity calc_ctrl
  end for;
end calc_ctrl_rtl_cfg;
